module nameduc (


);
endmodule
